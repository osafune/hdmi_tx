// c4e_pcmplay_core.v

// Generated using ACDS version 20.1 720

`timescale 1 ps / 1 ps
module c4e_pcmplay_core (
		output wire [11:0] bar_export,    //      bar.export
		input  wire        clk_100m_clk,  // clk_100m.clk
		input  wire        clk_25m_clk,   //  clk_25m.clk
		inout  wire [1:0]  gpio_export,   //     gpio.export
		input  wire        pcm_clk_128fs, //      pcm.clk_128fs
		output wire        pcm_fs,        //         .fs
		output wire [15:0] pcm_ldata,     //         .ldata
		output wire [15:0] pcm_rdata,     //         .rdata
		output wire        pcm_mute,      //         .mute
		input  wire        reset_reset_n, //    reset.reset_n
		output wire        sd_clk,        //       sd.clk
		output wire        sd_cmd,        //         .cmd
		input  wire        sd_dat0,       //         .dat0
		output wire        sd_dat3,       //         .dat3
		input  wire        sd_cd_n,       //         .cd_n
		output wire        sd_pwr,        //         .pwr
		output wire [12:0] sdr_addr,      //      sdr.addr
		output wire [1:0]  sdr_ba,        //         .ba
		output wire        sdr_cas_n,     //         .cas_n
		output wire        sdr_cke,       //         .cke
		output wire        sdr_cs_n,      //         .cs_n
		inout  wire [15:0] sdr_dq,        //         .dq
		output wire [1:0]  sdr_dqm,       //         .dqm
		output wire        sdr_ras_n,     //         .ras_n
		output wire        sdr_we_n,      //         .we_n
		input  wire        uart_rxd,      //     uart.rxd
		output wire        uart_txd,      //         .txd
		input  wire        vga_videoclk,  //      vga.videoclk
		output wire        vga_active,    //         .active
		output wire [7:0]  vga_rout,      //         .rout
		output wire [7:0]  vga_gout,      //         .gout
		output wire [7:0]  vga_bout,      //         .bout
		output wire        vga_hsync_n,   //         .hsync_n
		output wire        vga_vsync_n,   //         .vsync_n
		output wire        vga_csync_n    //         .csync_n
	);

	wire  [31:0] nios2_tiny_data_master_readdata;                          // mm_interconnect_0:nios2_tiny_data_master_readdata -> nios2_tiny:d_readdata
	wire         nios2_tiny_data_master_waitrequest;                       // mm_interconnect_0:nios2_tiny_data_master_waitrequest -> nios2_tiny:d_waitrequest
	wire         nios2_tiny_data_master_debugaccess;                       // nios2_tiny:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_tiny_data_master_debugaccess
	wire  [28:0] nios2_tiny_data_master_address;                           // nios2_tiny:d_address -> mm_interconnect_0:nios2_tiny_data_master_address
	wire   [3:0] nios2_tiny_data_master_byteenable;                        // nios2_tiny:d_byteenable -> mm_interconnect_0:nios2_tiny_data_master_byteenable
	wire         nios2_tiny_data_master_read;                              // nios2_tiny:d_read -> mm_interconnect_0:nios2_tiny_data_master_read
	wire         nios2_tiny_data_master_write;                             // nios2_tiny:d_write -> mm_interconnect_0:nios2_tiny_data_master_write
	wire  [31:0] nios2_tiny_data_master_writedata;                         // nios2_tiny:d_writedata -> mm_interconnect_0:nios2_tiny_data_master_writedata
	wire  [31:0] nios2_tiny_instruction_master_readdata;                   // mm_interconnect_0:nios2_tiny_instruction_master_readdata -> nios2_tiny:i_readdata
	wire         nios2_tiny_instruction_master_waitrequest;                // mm_interconnect_0:nios2_tiny_instruction_master_waitrequest -> nios2_tiny:i_waitrequest
	wire  [27:0] nios2_tiny_instruction_master_address;                    // nios2_tiny:i_address -> mm_interconnect_0:nios2_tiny_instruction_master_address
	wire         nios2_tiny_instruction_master_read;                       // nios2_tiny:i_read -> mm_interconnect_0:nios2_tiny_instruction_master_read
	wire         vga_m1_waitrequest;                                       // mm_interconnect_0:vga_m1_waitrequest -> vga:avm_m1_waitrequest
	wire  [31:0] vga_m1_readdata;                                          // mm_interconnect_0:vga_m1_readdata -> vga:avm_m1_readdata
	wire  [31:0] vga_m1_address;                                           // vga:avm_m1_address -> mm_interconnect_0:vga_m1_address
	wire         vga_m1_read;                                              // vga:avm_m1_read -> mm_interconnect_0:vga_m1_read
	wire         vga_m1_readdatavalid;                                     // mm_interconnect_0:vga_m1_readdatavalid -> vga:avm_m1_readdatavalid
	wire   [8:0] vga_m1_burstcount;                                        // vga:avm_m1_burstcount -> mm_interconnect_0:vga_m1_burstcount
	wire  [31:0] mm_interconnect_0_nios2_tiny_debug_mem_slave_readdata;    // nios2_tiny:debug_mem_slave_readdata -> mm_interconnect_0:nios2_tiny_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_tiny_debug_mem_slave_waitrequest; // nios2_tiny:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_tiny_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_tiny_debug_mem_slave_debugaccess; // mm_interconnect_0:nios2_tiny_debug_mem_slave_debugaccess -> nios2_tiny:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_tiny_debug_mem_slave_address;     // mm_interconnect_0:nios2_tiny_debug_mem_slave_address -> nios2_tiny:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_tiny_debug_mem_slave_read;        // mm_interconnect_0:nios2_tiny_debug_mem_slave_read -> nios2_tiny:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_tiny_debug_mem_slave_byteenable;  // mm_interconnect_0:nios2_tiny_debug_mem_slave_byteenable -> nios2_tiny:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_tiny_debug_mem_slave_write;       // mm_interconnect_0:nios2_tiny_debug_mem_slave_write -> nios2_tiny:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_tiny_debug_mem_slave_writedata;   // mm_interconnect_0:nios2_tiny_debug_mem_slave_writedata -> nios2_tiny:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_peripheral_bridge_s0_readdata;          // peripheral_bridge:s0_readdata -> mm_interconnect_0:peripheral_bridge_s0_readdata
	wire         mm_interconnect_0_peripheral_bridge_s0_waitrequest;       // peripheral_bridge:s0_waitrequest -> mm_interconnect_0:peripheral_bridge_s0_waitrequest
	wire         mm_interconnect_0_peripheral_bridge_s0_debugaccess;       // mm_interconnect_0:peripheral_bridge_s0_debugaccess -> peripheral_bridge:s0_debugaccess
	wire   [8:0] mm_interconnect_0_peripheral_bridge_s0_address;           // mm_interconnect_0:peripheral_bridge_s0_address -> peripheral_bridge:s0_address
	wire         mm_interconnect_0_peripheral_bridge_s0_read;              // mm_interconnect_0:peripheral_bridge_s0_read -> peripheral_bridge:s0_read
	wire   [3:0] mm_interconnect_0_peripheral_bridge_s0_byteenable;        // mm_interconnect_0:peripheral_bridge_s0_byteenable -> peripheral_bridge:s0_byteenable
	wire         mm_interconnect_0_peripheral_bridge_s0_readdatavalid;     // peripheral_bridge:s0_readdatavalid -> mm_interconnect_0:peripheral_bridge_s0_readdatavalid
	wire         mm_interconnect_0_peripheral_bridge_s0_write;             // mm_interconnect_0:peripheral_bridge_s0_write -> peripheral_bridge:s0_write
	wire  [31:0] mm_interconnect_0_peripheral_bridge_s0_writedata;         // mm_interconnect_0:peripheral_bridge_s0_writedata -> peripheral_bridge:s0_writedata
	wire   [0:0] mm_interconnect_0_peripheral_bridge_s0_burstcount;        // mm_interconnect_0:peripheral_bridge_s0_burstcount -> peripheral_bridge:s0_burstcount
	wire  [31:0] mm_interconnect_0_pcm_s0_readdata;                        // pcm:avs_readdata -> mm_interconnect_0:pcm_s0_readdata
	wire   [1:0] mm_interconnect_0_pcm_s0_address;                         // mm_interconnect_0:pcm_s0_address -> pcm:avs_address
	wire         mm_interconnect_0_pcm_s0_read;                            // mm_interconnect_0:pcm_s0_read -> pcm:avs_read
	wire         mm_interconnect_0_pcm_s0_write;                           // mm_interconnect_0:pcm_s0_write -> pcm:avs_write
	wire  [31:0] mm_interconnect_0_pcm_s0_writedata;                       // mm_interconnect_0:pcm_s0_writedata -> pcm:avs_writedata
	wire         mm_interconnect_0_sdram_s1_chipselect;                    // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;                      // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                   // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [23:0] mm_interconnect_0_sdram_s1_address;                       // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                          // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;                    // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                 // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                         // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;                     // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire         mm_interconnect_0_boot_s1_chipselect;                     // mm_interconnect_0:boot_s1_chipselect -> boot:chipselect
	wire  [31:0] mm_interconnect_0_boot_s1_readdata;                       // boot:readdata -> mm_interconnect_0:boot_s1_readdata
	wire  [11:0] mm_interconnect_0_boot_s1_address;                        // mm_interconnect_0:boot_s1_address -> boot:address
	wire   [3:0] mm_interconnect_0_boot_s1_byteenable;                     // mm_interconnect_0:boot_s1_byteenable -> boot:byteenable
	wire         mm_interconnect_0_boot_s1_write;                          // mm_interconnect_0:boot_s1_write -> boot:write
	wire  [31:0] mm_interconnect_0_boot_s1_writedata;                      // mm_interconnect_0:boot_s1_writedata -> boot:writedata
	wire         mm_interconnect_0_boot_s1_clken;                          // mm_interconnect_0:boot_s1_clken -> boot:clken
	wire  [31:0] mm_interconnect_0_peridot_sdif_0_s1_readdata;             // peridot_sdif_0:avs_readdata -> mm_interconnect_0:peridot_sdif_0_s1_readdata
	wire   [1:0] mm_interconnect_0_peridot_sdif_0_s1_address;              // mm_interconnect_0:peridot_sdif_0_s1_address -> peridot_sdif_0:avs_address
	wire         mm_interconnect_0_peridot_sdif_0_s1_read;                 // mm_interconnect_0:peridot_sdif_0_s1_read -> peridot_sdif_0:avs_read
	wire         mm_interconnect_0_peridot_sdif_0_s1_write;                // mm_interconnect_0:peridot_sdif_0_s1_write -> peridot_sdif_0:avs_write
	wire  [31:0] mm_interconnect_0_peridot_sdif_0_s1_writedata;            // mm_interconnect_0:peridot_sdif_0_s1_writedata -> peridot_sdif_0:avs_writedata
	wire         peripheral_bridge_m0_waitrequest;                         // mm_interconnect_1:peripheral_bridge_m0_waitrequest -> peripheral_bridge:m0_waitrequest
	wire  [31:0] peripheral_bridge_m0_readdata;                            // mm_interconnect_1:peripheral_bridge_m0_readdata -> peripheral_bridge:m0_readdata
	wire         peripheral_bridge_m0_debugaccess;                         // peripheral_bridge:m0_debugaccess -> mm_interconnect_1:peripheral_bridge_m0_debugaccess
	wire   [8:0] peripheral_bridge_m0_address;                             // peripheral_bridge:m0_address -> mm_interconnect_1:peripheral_bridge_m0_address
	wire         peripheral_bridge_m0_read;                                // peripheral_bridge:m0_read -> mm_interconnect_1:peripheral_bridge_m0_read
	wire   [3:0] peripheral_bridge_m0_byteenable;                          // peripheral_bridge:m0_byteenable -> mm_interconnect_1:peripheral_bridge_m0_byteenable
	wire         peripheral_bridge_m0_readdatavalid;                       // mm_interconnect_1:peripheral_bridge_m0_readdatavalid -> peripheral_bridge:m0_readdatavalid
	wire  [31:0] peripheral_bridge_m0_writedata;                           // peripheral_bridge:m0_writedata -> mm_interconnect_1:peripheral_bridge_m0_writedata
	wire         peripheral_bridge_m0_write;                               // peripheral_bridge:m0_write -> mm_interconnect_1:peripheral_bridge_m0_write
	wire   [0:0] peripheral_bridge_m0_burstcount;                          // peripheral_bridge:m0_burstcount -> mm_interconnect_1:peripheral_bridge_m0_burstcount
	wire  [31:0] mm_interconnect_1_sysid_control_slave_readdata;           // sysid:readdata -> mm_interconnect_1:sysid_control_slave_readdata
	wire   [0:0] mm_interconnect_1_sysid_control_slave_address;            // mm_interconnect_1:sysid_control_slave_address -> sysid:address
	wire  [31:0] mm_interconnect_1_vga_csr_readdata;                       // vga:avs_csr_readdata -> mm_interconnect_1:vga_csr_readdata
	wire   [1:0] mm_interconnect_1_vga_csr_address;                        // mm_interconnect_1:vga_csr_address -> vga:avs_csr_address
	wire         mm_interconnect_1_vga_csr_read;                           // mm_interconnect_1:vga_csr_read -> vga:avs_csr_read
	wire         mm_interconnect_1_vga_csr_write;                          // mm_interconnect_1:vga_csr_write -> vga:avs_csr_write
	wire  [31:0] mm_interconnect_1_vga_csr_writedata;                      // mm_interconnect_1:vga_csr_writedata -> vga:avs_csr_writedata
	wire         mm_interconnect_1_systimer_s1_chipselect;                 // mm_interconnect_1:systimer_s1_chipselect -> systimer:chipselect
	wire  [15:0] mm_interconnect_1_systimer_s1_readdata;                   // systimer:readdata -> mm_interconnect_1:systimer_s1_readdata
	wire   [2:0] mm_interconnect_1_systimer_s1_address;                    // mm_interconnect_1:systimer_s1_address -> systimer:address
	wire         mm_interconnect_1_systimer_s1_write;                      // mm_interconnect_1:systimer_s1_write -> systimer:write_n
	wire  [15:0] mm_interconnect_1_systimer_s1_writedata;                  // mm_interconnect_1:systimer_s1_writedata -> systimer:writedata
	wire         mm_interconnect_1_gpio_s1_chipselect;                     // mm_interconnect_1:gpio_s1_chipselect -> gpio:chipselect
	wire  [31:0] mm_interconnect_1_gpio_s1_readdata;                       // gpio:readdata -> mm_interconnect_1:gpio_s1_readdata
	wire   [1:0] mm_interconnect_1_gpio_s1_address;                        // mm_interconnect_1:gpio_s1_address -> gpio:address
	wire         mm_interconnect_1_gpio_s1_write;                          // mm_interconnect_1:gpio_s1_write -> gpio:write_n
	wire  [31:0] mm_interconnect_1_gpio_s1_writedata;                      // mm_interconnect_1:gpio_s1_writedata -> gpio:writedata
	wire         mm_interconnect_1_sysuart_s1_chipselect;                  // mm_interconnect_1:sysuart_s1_chipselect -> sysuart:chipselect
	wire  [15:0] mm_interconnect_1_sysuart_s1_readdata;                    // sysuart:readdata -> mm_interconnect_1:sysuart_s1_readdata
	wire   [2:0] mm_interconnect_1_sysuart_s1_address;                     // mm_interconnect_1:sysuart_s1_address -> sysuart:address
	wire         mm_interconnect_1_sysuart_s1_read;                        // mm_interconnect_1:sysuart_s1_read -> sysuart:read_n
	wire         mm_interconnect_1_sysuart_s1_begintransfer;               // mm_interconnect_1:sysuart_s1_begintransfer -> sysuart:begintransfer
	wire         mm_interconnect_1_sysuart_s1_write;                       // mm_interconnect_1:sysuart_s1_write -> sysuart:write_n
	wire  [15:0] mm_interconnect_1_sysuart_s1_writedata;                   // mm_interconnect_1:sysuart_s1_writedata -> sysuart:writedata
	wire         mm_interconnect_1_barcolor_s1_chipselect;                 // mm_interconnect_1:barcolor_s1_chipselect -> barcolor:chipselect
	wire  [31:0] mm_interconnect_1_barcolor_s1_readdata;                   // barcolor:readdata -> mm_interconnect_1:barcolor_s1_readdata
	wire   [1:0] mm_interconnect_1_barcolor_s1_address;                    // mm_interconnect_1:barcolor_s1_address -> barcolor:address
	wire         mm_interconnect_1_barcolor_s1_write;                      // mm_interconnect_1:barcolor_s1_write -> barcolor:write_n
	wire  [31:0] mm_interconnect_1_barcolor_s1_writedata;                  // mm_interconnect_1:barcolor_s1_writedata -> barcolor:writedata
	wire         irq_mapper_receiver1_irq;                                 // peridot_sdif_0:ins_irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver4_irq;                                 // pcm:ins_irq -> irq_mapper:receiver4_irq
	wire  [31:0] nios2_tiny_irq_irq;                                       // irq_mapper:sender_irq -> nios2_tiny:irq
	wire         irq_mapper_receiver0_irq;                                 // irq_synchronizer:sender_irq -> irq_mapper:receiver0_irq
	wire   [0:0] irq_synchronizer_receiver_irq;                            // systimer:irq -> irq_synchronizer:receiver_irq
	wire         irq_mapper_receiver2_irq;                                 // irq_synchronizer_001:sender_irq -> irq_mapper:receiver2_irq
	wire   [0:0] irq_synchronizer_001_receiver_irq;                        // sysuart:irq -> irq_synchronizer_001:receiver_irq
	wire         irq_mapper_receiver3_irq;                                 // irq_synchronizer_002:sender_irq -> irq_mapper:receiver3_irq
	wire   [0:0] irq_synchronizer_002_receiver_irq;                        // vga:ins_csr_irq -> irq_synchronizer_002:receiver_irq
	wire         rst_controller_reset_out_reset;                           // rst_controller:reset_out -> [barcolor:reset_n, gpio:reset_n, irq_synchronizer:receiver_reset, irq_synchronizer_001:receiver_reset, irq_synchronizer_002:receiver_reset, mm_interconnect_0:peripheral_bridge_reset_reset_bridge_in_reset_reset, mm_interconnect_1:peripheral_bridge_reset_reset_bridge_in_reset_reset, peripheral_bridge:reset, sysid:reset_n, systimer:reset_n, sysuart:reset_n, vga:csi_csr_reset]
	wire         rst_controller_001_reset_out_reset;                       // rst_controller_001:reset_out -> [boot:reset, irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, irq_synchronizer_002:sender_reset, mm_interconnect_0:nios2_tiny_reset_reset_bridge_in_reset_reset, nios2_tiny:reset_n, rst_translator:in_reset]
	wire         rst_controller_001_reset_out_reset_req;                   // rst_controller_001:reset_req -> [boot:reset_req, nios2_tiny:reset_req, rst_translator:reset_req_in]
	wire         nios2_tiny_debug_reset_request_reset;                     // nios2_tiny:debug_reset_request -> rst_controller_001:reset_in1
	wire         rst_controller_002_reset_out_reset;                       // rst_controller_002:reset_out -> [mm_interconnect_0:pcm_reset_reset_bridge_in_reset_reset, pcm:csi_reset, peridot_sdif_0:csi_reset, sdram:reset_n]
	wire         rst_controller_003_reset_out_reset;                       // rst_controller_003:reset_out -> mm_interconnect_0:vga_reset_reset_bridge_in_reset_reset

	c4e_pcmplay_core_barcolor barcolor (
		.clk        (clk_25m_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_1_barcolor_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_barcolor_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_barcolor_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_barcolor_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_barcolor_s1_readdata),   //                    .readdata
		.out_port   (bar_export)                                // external_connection.export
	);

	c4e_pcmplay_core_boot boot (
		.clk        (clk_100m_clk),                           //   clk1.clk
		.address    (mm_interconnect_0_boot_s1_address),      //     s1.address
		.clken      (mm_interconnect_0_boot_s1_clken),        //       .clken
		.chipselect (mm_interconnect_0_boot_s1_chipselect),   //       .chipselect
		.write      (mm_interconnect_0_boot_s1_write),        //       .write
		.readdata   (mm_interconnect_0_boot_s1_readdata),     //       .readdata
		.writedata  (mm_interconnect_0_boot_s1_writedata),    //       .writedata
		.byteenable (mm_interconnect_0_boot_s1_byteenable),   //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),     // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req), //       .reset_req
		.freeze     (1'b0)                                    // (terminated)
	);

	c4e_pcmplay_core_gpio gpio (
		.clk        (clk_25m_clk),                          //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_1_gpio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_gpio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_gpio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_gpio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_gpio_s1_readdata),   //                    .readdata
		.bidir_port (gpio_export)                           // external_connection.export
	);

	c4e_pcmplay_core_nios2_tiny nios2_tiny (
		.clk                                 (clk_100m_clk),                                             //                       clk.clk
		.reset_n                             (~rst_controller_001_reset_out_reset),                      //                     reset.reset_n
		.reset_req                           (rst_controller_001_reset_out_reset_req),                   //                          .reset_req
		.d_address                           (nios2_tiny_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_tiny_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_tiny_data_master_read),                              //                          .read
		.d_readdata                          (nios2_tiny_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_tiny_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_tiny_data_master_write),                             //                          .write
		.d_writedata                         (nios2_tiny_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_tiny_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_tiny_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_tiny_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_tiny_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_tiny_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_tiny_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_tiny_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_tiny_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_tiny_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_tiny_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_tiny_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_tiny_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_tiny_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_tiny_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_tiny_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                          // custom_instruction_master.readra
	);

	pcm_component pcm (
		.csi_clk       (clk_100m_clk),                       //  clock.clk
		.csi_reset     (rst_controller_002_reset_out_reset), //  reset.reset
		.avs_address   (mm_interconnect_0_pcm_s0_address),   //     s0.address
		.avs_read      (mm_interconnect_0_pcm_s0_read),      //       .read
		.avs_readdata  (mm_interconnect_0_pcm_s0_readdata),  //       .readdata
		.avs_write     (mm_interconnect_0_pcm_s0_write),     //       .write
		.avs_writedata (mm_interconnect_0_pcm_s0_writedata), //       .writedata
		.ins_irq       (irq_mapper_receiver4_irq),           //    irs.irq
		.coe_128fs_clk (pcm_clk_128fs),                      // export.clk_128fs
		.coe_pcm_fs    (pcm_fs),                             //       .fs
		.coe_pcm_l     (pcm_ldata),                          //       .ldata
		.coe_pcm_r     (pcm_rdata),                          //       .rdata
		.coe_mute      (pcm_mute)                            //       .mute
	);

	peridot_sdif peridot_sdif_0 (
		.csi_clk       (clk_100m_clk),                                  //  clock.clk
		.csi_reset     (rst_controller_002_reset_out_reset),            //  reset.reset
		.avs_address   (mm_interconnect_0_peridot_sdif_0_s1_address),   //     s1.address
		.avs_read      (mm_interconnect_0_peridot_sdif_0_s1_read),      //       .read
		.avs_readdata  (mm_interconnect_0_peridot_sdif_0_s1_readdata),  //       .readdata
		.avs_write     (mm_interconnect_0_peridot_sdif_0_s1_write),     //       .write
		.avs_writedata (mm_interconnect_0_peridot_sdif_0_s1_writedata), //       .writedata
		.ins_irq       (irq_mapper_receiver1_irq),                      //    irq.irq
		.coe_sd_clk    (sd_clk),                                        // export.clk
		.coe_sd_cmd    (sd_cmd),                                        //       .cmd
		.coe_sd_dat0   (sd_dat0),                                       //       .dat0
		.coe_sd_dat3   (sd_dat3),                                       //       .dat3
		.coe_sd_cd_n   (sd_cd_n),                                       //       .cd_n
		.coe_sd_pwr    (sd_pwr)                                         //       .pwr
	);

	altera_avalon_mm_bridge #(
		.DATA_WIDTH        (32),
		.SYMBOL_WIDTH      (8),
		.HDL_ADDR_WIDTH    (9),
		.BURSTCOUNT_WIDTH  (1),
		.PIPELINE_COMMAND  (1),
		.PIPELINE_RESPONSE (1)
	) peripheral_bridge (
		.clk              (clk_25m_clk),                                          //   clk.clk
		.reset            (rst_controller_reset_out_reset),                       // reset.reset
		.s0_waitrequest   (mm_interconnect_0_peripheral_bridge_s0_waitrequest),   //    s0.waitrequest
		.s0_readdata      (mm_interconnect_0_peripheral_bridge_s0_readdata),      //      .readdata
		.s0_readdatavalid (mm_interconnect_0_peripheral_bridge_s0_readdatavalid), //      .readdatavalid
		.s0_burstcount    (mm_interconnect_0_peripheral_bridge_s0_burstcount),    //      .burstcount
		.s0_writedata     (mm_interconnect_0_peripheral_bridge_s0_writedata),     //      .writedata
		.s0_address       (mm_interconnect_0_peripheral_bridge_s0_address),       //      .address
		.s0_write         (mm_interconnect_0_peripheral_bridge_s0_write),         //      .write
		.s0_read          (mm_interconnect_0_peripheral_bridge_s0_read),          //      .read
		.s0_byteenable    (mm_interconnect_0_peripheral_bridge_s0_byteenable),    //      .byteenable
		.s0_debugaccess   (mm_interconnect_0_peripheral_bridge_s0_debugaccess),   //      .debugaccess
		.m0_waitrequest   (peripheral_bridge_m0_waitrequest),                     //    m0.waitrequest
		.m0_readdata      (peripheral_bridge_m0_readdata),                        //      .readdata
		.m0_readdatavalid (peripheral_bridge_m0_readdatavalid),                   //      .readdatavalid
		.m0_burstcount    (peripheral_bridge_m0_burstcount),                      //      .burstcount
		.m0_writedata     (peripheral_bridge_m0_writedata),                       //      .writedata
		.m0_address       (peripheral_bridge_m0_address),                         //      .address
		.m0_write         (peripheral_bridge_m0_write),                           //      .write
		.m0_read          (peripheral_bridge_m0_read),                            //      .read
		.m0_byteenable    (peripheral_bridge_m0_byteenable),                      //      .byteenable
		.m0_debugaccess   (peripheral_bridge_m0_debugaccess),                     //      .debugaccess
		.s0_response      (),                                                     // (terminated)
		.m0_response      (2'b00)                                                 // (terminated)
	);

	c4e_pcmplay_core_sdram sdram (
		.clk            (clk_100m_clk),                             //   clk.clk
		.reset_n        (~rst_controller_002_reset_out_reset),      // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdr_addr),                                 //  wire.export
		.zs_ba          (sdr_ba),                                   //      .export
		.zs_cas_n       (sdr_cas_n),                                //      .export
		.zs_cke         (sdr_cke),                                  //      .export
		.zs_cs_n        (sdr_cs_n),                                 //      .export
		.zs_dq          (sdr_dq),                                   //      .export
		.zs_dqm         (sdr_dqm),                                  //      .export
		.zs_ras_n       (sdr_ras_n),                                //      .export
		.zs_we_n        (sdr_we_n)                                  //      .export
	);

	c4e_pcmplay_core_sysid sysid (
		.clock    (clk_25m_clk),                                    //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //         reset.reset_n
		.readdata (mm_interconnect_1_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_1_sysid_control_slave_address)   //              .address
	);

	c4e_pcmplay_core_systimer systimer (
		.clk        (clk_25m_clk),                              //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          // reset.reset_n
		.address    (mm_interconnect_1_systimer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_1_systimer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_1_systimer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_1_systimer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_1_systimer_s1_write),     //      .write_n
		.irq        (irq_synchronizer_receiver_irq)             //   irq.irq
	);

	c4e_pcmplay_core_sysuart sysuart (
		.clk           (clk_25m_clk),                                //                 clk.clk
		.reset_n       (~rst_controller_reset_out_reset),            //               reset.reset_n
		.address       (mm_interconnect_1_sysuart_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_1_sysuart_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_1_sysuart_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_1_sysuart_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_1_sysuart_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_1_sysuart_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_1_sysuart_s1_readdata),      //                    .readdata
		.rxd           (uart_rxd),                                   // external_connection.export
		.txd           (uart_txd),                                   //                    .export
		.irq           (irq_synchronizer_001_receiver_irq)           //                 irq.irq
	);

	peridot_vga #(
		.DEVICE_FAMILY       ("Cyclone IV E"),
		.FIFORESETCOUNT      (9),
		.FIFODEPTH_WIDTH     (10),
		.VIDEO_INTERFACE     ("PARALLEL"),
		.VGACLOCK_FREQUENCY  (74250000),
		.H_TOTAL             (1650),
		.H_SYNC              (40),
		.H_BACKP             (220),
		.H_ACTIVE            (1280),
		.V_TOTAL             (750),
		.V_SYNC              (5),
		.V_BACKP             (20),
		.V_ACTIVE            (720),
		.USE_AUDIOSTREAM     ("OFF"),
		.BURSTCOUNT_WIDTH    (8),
		.LINEOFFSETBYTES     (2560),
		.PIXEL_DATAORDER     ("BYTE"),
		.PIXEL_COLORORDER    ("RGB565"),
		.PCMSAMPLE_FREQUENCY (44100)
	) vga (
		.csi_csr_clk          (clk_25m_clk),                         // csr_clk.clk
		.csi_csr_reset        (rst_controller_reset_out_reset),      //   reset.reset
		.avs_csr_address      (mm_interconnect_1_vga_csr_address),   //     csr.address
		.avs_csr_read         (mm_interconnect_1_vga_csr_read),      //        .read
		.avs_csr_readdata     (mm_interconnect_1_vga_csr_readdata),  //        .readdata
		.avs_csr_write        (mm_interconnect_1_vga_csr_write),     //        .write
		.avs_csr_writedata    (mm_interconnect_1_vga_csr_writedata), //        .writedata
		.ins_csr_irq          (irq_synchronizer_002_receiver_irq),   // irq_csr.irq
		.csi_m1_clk           (clk_100m_clk),                        //  m1_clk.clk
		.avm_m1_waitrequest   (vga_m1_waitrequest),                  //      m1.waitrequest
		.avm_m1_address       (vga_m1_address),                      //        .address
		.avm_m1_read          (vga_m1_read),                         //        .read
		.avm_m1_readdata      (vga_m1_readdata),                     //        .readdata
		.avm_m1_readdatavalid (vga_m1_readdatavalid),                //        .readdatavalid
		.avm_m1_burstcount    (vga_m1_burstcount),                   //        .burstcount
		.coe_vga_clk          (vga_videoclk),                        //     vga.videoclk
		.coe_vga_active       (vga_active),                          //        .active
		.coe_vga_rout         (vga_rout),                            //        .rout
		.coe_vga_gout         (vga_gout),                            //        .gout
		.coe_vga_bout         (vga_bout),                            //        .bout
		.coe_vga_hsync_n      (vga_hsync_n),                         //        .hsync_n
		.coe_vga_vsync_n      (vga_vsync_n),                         //        .vsync_n
		.coe_vga_csync_n      (vga_csync_n),                         //        .csync_n
		.coe_pcm_fs           (1'b0),                                // (terminated)
		.coe_pcm_l            (24'b000000000000000000000000),        // (terminated)
		.coe_pcm_r            (24'b000000000000000000000000),        // (terminated)
		.coe_ser_clk          (1'b0),                                // (terminated)
		.coe_ser_x5clk        (1'b0),                                // (terminated)
		.coe_ser_data         (),                                    // (terminated)
		.coe_ser_data_n       (),                                    // (terminated)
		.coe_ser_clock        (),                                    // (terminated)
		.coe_ser_clock_n      ()                                     // (terminated)
	);

	c4e_pcmplay_core_mm_interconnect_0 mm_interconnect_0 (
		.core_clk_clk_clk                                    (clk_100m_clk),                                             //                                  core_clk_clk.clk
		.peri_clk_clk_clk                                    (clk_25m_clk),                                              //                                  peri_clk_clk.clk
		.nios2_tiny_reset_reset_bridge_in_reset_reset        (rst_controller_001_reset_out_reset),                       //        nios2_tiny_reset_reset_bridge_in_reset.reset
		.pcm_reset_reset_bridge_in_reset_reset               (rst_controller_002_reset_out_reset),                       //               pcm_reset_reset_bridge_in_reset.reset
		.peripheral_bridge_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                           // peripheral_bridge_reset_reset_bridge_in_reset.reset
		.vga_reset_reset_bridge_in_reset_reset               (rst_controller_003_reset_out_reset),                       //               vga_reset_reset_bridge_in_reset.reset
		.nios2_tiny_data_master_address                      (nios2_tiny_data_master_address),                           //                        nios2_tiny_data_master.address
		.nios2_tiny_data_master_waitrequest                  (nios2_tiny_data_master_waitrequest),                       //                                              .waitrequest
		.nios2_tiny_data_master_byteenable                   (nios2_tiny_data_master_byteenable),                        //                                              .byteenable
		.nios2_tiny_data_master_read                         (nios2_tiny_data_master_read),                              //                                              .read
		.nios2_tiny_data_master_readdata                     (nios2_tiny_data_master_readdata),                          //                                              .readdata
		.nios2_tiny_data_master_write                        (nios2_tiny_data_master_write),                             //                                              .write
		.nios2_tiny_data_master_writedata                    (nios2_tiny_data_master_writedata),                         //                                              .writedata
		.nios2_tiny_data_master_debugaccess                  (nios2_tiny_data_master_debugaccess),                       //                                              .debugaccess
		.nios2_tiny_instruction_master_address               (nios2_tiny_instruction_master_address),                    //                 nios2_tiny_instruction_master.address
		.nios2_tiny_instruction_master_waitrequest           (nios2_tiny_instruction_master_waitrequest),                //                                              .waitrequest
		.nios2_tiny_instruction_master_read                  (nios2_tiny_instruction_master_read),                       //                                              .read
		.nios2_tiny_instruction_master_readdata              (nios2_tiny_instruction_master_readdata),                   //                                              .readdata
		.vga_m1_address                                      (vga_m1_address),                                           //                                        vga_m1.address
		.vga_m1_waitrequest                                  (vga_m1_waitrequest),                                       //                                              .waitrequest
		.vga_m1_burstcount                                   (vga_m1_burstcount),                                        //                                              .burstcount
		.vga_m1_read                                         (vga_m1_read),                                              //                                              .read
		.vga_m1_readdata                                     (vga_m1_readdata),                                          //                                              .readdata
		.vga_m1_readdatavalid                                (vga_m1_readdatavalid),                                     //                                              .readdatavalid
		.boot_s1_address                                     (mm_interconnect_0_boot_s1_address),                        //                                       boot_s1.address
		.boot_s1_write                                       (mm_interconnect_0_boot_s1_write),                          //                                              .write
		.boot_s1_readdata                                    (mm_interconnect_0_boot_s1_readdata),                       //                                              .readdata
		.boot_s1_writedata                                   (mm_interconnect_0_boot_s1_writedata),                      //                                              .writedata
		.boot_s1_byteenable                                  (mm_interconnect_0_boot_s1_byteenable),                     //                                              .byteenable
		.boot_s1_chipselect                                  (mm_interconnect_0_boot_s1_chipselect),                     //                                              .chipselect
		.boot_s1_clken                                       (mm_interconnect_0_boot_s1_clken),                          //                                              .clken
		.nios2_tiny_debug_mem_slave_address                  (mm_interconnect_0_nios2_tiny_debug_mem_slave_address),     //                    nios2_tiny_debug_mem_slave.address
		.nios2_tiny_debug_mem_slave_write                    (mm_interconnect_0_nios2_tiny_debug_mem_slave_write),       //                                              .write
		.nios2_tiny_debug_mem_slave_read                     (mm_interconnect_0_nios2_tiny_debug_mem_slave_read),        //                                              .read
		.nios2_tiny_debug_mem_slave_readdata                 (mm_interconnect_0_nios2_tiny_debug_mem_slave_readdata),    //                                              .readdata
		.nios2_tiny_debug_mem_slave_writedata                (mm_interconnect_0_nios2_tiny_debug_mem_slave_writedata),   //                                              .writedata
		.nios2_tiny_debug_mem_slave_byteenable               (mm_interconnect_0_nios2_tiny_debug_mem_slave_byteenable),  //                                              .byteenable
		.nios2_tiny_debug_mem_slave_waitrequest              (mm_interconnect_0_nios2_tiny_debug_mem_slave_waitrequest), //                                              .waitrequest
		.nios2_tiny_debug_mem_slave_debugaccess              (mm_interconnect_0_nios2_tiny_debug_mem_slave_debugaccess), //                                              .debugaccess
		.pcm_s0_address                                      (mm_interconnect_0_pcm_s0_address),                         //                                        pcm_s0.address
		.pcm_s0_write                                        (mm_interconnect_0_pcm_s0_write),                           //                                              .write
		.pcm_s0_read                                         (mm_interconnect_0_pcm_s0_read),                            //                                              .read
		.pcm_s0_readdata                                     (mm_interconnect_0_pcm_s0_readdata),                        //                                              .readdata
		.pcm_s0_writedata                                    (mm_interconnect_0_pcm_s0_writedata),                       //                                              .writedata
		.peridot_sdif_0_s1_address                           (mm_interconnect_0_peridot_sdif_0_s1_address),              //                             peridot_sdif_0_s1.address
		.peridot_sdif_0_s1_write                             (mm_interconnect_0_peridot_sdif_0_s1_write),                //                                              .write
		.peridot_sdif_0_s1_read                              (mm_interconnect_0_peridot_sdif_0_s1_read),                 //                                              .read
		.peridot_sdif_0_s1_readdata                          (mm_interconnect_0_peridot_sdif_0_s1_readdata),             //                                              .readdata
		.peridot_sdif_0_s1_writedata                         (mm_interconnect_0_peridot_sdif_0_s1_writedata),            //                                              .writedata
		.peripheral_bridge_s0_address                        (mm_interconnect_0_peripheral_bridge_s0_address),           //                          peripheral_bridge_s0.address
		.peripheral_bridge_s0_write                          (mm_interconnect_0_peripheral_bridge_s0_write),             //                                              .write
		.peripheral_bridge_s0_read                           (mm_interconnect_0_peripheral_bridge_s0_read),              //                                              .read
		.peripheral_bridge_s0_readdata                       (mm_interconnect_0_peripheral_bridge_s0_readdata),          //                                              .readdata
		.peripheral_bridge_s0_writedata                      (mm_interconnect_0_peripheral_bridge_s0_writedata),         //                                              .writedata
		.peripheral_bridge_s0_burstcount                     (mm_interconnect_0_peripheral_bridge_s0_burstcount),        //                                              .burstcount
		.peripheral_bridge_s0_byteenable                     (mm_interconnect_0_peripheral_bridge_s0_byteenable),        //                                              .byteenable
		.peripheral_bridge_s0_readdatavalid                  (mm_interconnect_0_peripheral_bridge_s0_readdatavalid),     //                                              .readdatavalid
		.peripheral_bridge_s0_waitrequest                    (mm_interconnect_0_peripheral_bridge_s0_waitrequest),       //                                              .waitrequest
		.peripheral_bridge_s0_debugaccess                    (mm_interconnect_0_peripheral_bridge_s0_debugaccess),       //                                              .debugaccess
		.sdram_s1_address                                    (mm_interconnect_0_sdram_s1_address),                       //                                      sdram_s1.address
		.sdram_s1_write                                      (mm_interconnect_0_sdram_s1_write),                         //                                              .write
		.sdram_s1_read                                       (mm_interconnect_0_sdram_s1_read),                          //                                              .read
		.sdram_s1_readdata                                   (mm_interconnect_0_sdram_s1_readdata),                      //                                              .readdata
		.sdram_s1_writedata                                  (mm_interconnect_0_sdram_s1_writedata),                     //                                              .writedata
		.sdram_s1_byteenable                                 (mm_interconnect_0_sdram_s1_byteenable),                    //                                              .byteenable
		.sdram_s1_readdatavalid                              (mm_interconnect_0_sdram_s1_readdatavalid),                 //                                              .readdatavalid
		.sdram_s1_waitrequest                                (mm_interconnect_0_sdram_s1_waitrequest),                   //                                              .waitrequest
		.sdram_s1_chipselect                                 (mm_interconnect_0_sdram_s1_chipselect)                     //                                              .chipselect
	);

	c4e_pcmplay_core_mm_interconnect_1 mm_interconnect_1 (
		.peri_clk_clk_clk                                    (clk_25m_clk),                                    //                                  peri_clk_clk.clk
		.peripheral_bridge_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                 // peripheral_bridge_reset_reset_bridge_in_reset.reset
		.peripheral_bridge_m0_address                        (peripheral_bridge_m0_address),                   //                          peripheral_bridge_m0.address
		.peripheral_bridge_m0_waitrequest                    (peripheral_bridge_m0_waitrequest),               //                                              .waitrequest
		.peripheral_bridge_m0_burstcount                     (peripheral_bridge_m0_burstcount),                //                                              .burstcount
		.peripheral_bridge_m0_byteenable                     (peripheral_bridge_m0_byteenable),                //                                              .byteenable
		.peripheral_bridge_m0_read                           (peripheral_bridge_m0_read),                      //                                              .read
		.peripheral_bridge_m0_readdata                       (peripheral_bridge_m0_readdata),                  //                                              .readdata
		.peripheral_bridge_m0_readdatavalid                  (peripheral_bridge_m0_readdatavalid),             //                                              .readdatavalid
		.peripheral_bridge_m0_write                          (peripheral_bridge_m0_write),                     //                                              .write
		.peripheral_bridge_m0_writedata                      (peripheral_bridge_m0_writedata),                 //                                              .writedata
		.peripheral_bridge_m0_debugaccess                    (peripheral_bridge_m0_debugaccess),               //                                              .debugaccess
		.barcolor_s1_address                                 (mm_interconnect_1_barcolor_s1_address),          //                                   barcolor_s1.address
		.barcolor_s1_write                                   (mm_interconnect_1_barcolor_s1_write),            //                                              .write
		.barcolor_s1_readdata                                (mm_interconnect_1_barcolor_s1_readdata),         //                                              .readdata
		.barcolor_s1_writedata                               (mm_interconnect_1_barcolor_s1_writedata),        //                                              .writedata
		.barcolor_s1_chipselect                              (mm_interconnect_1_barcolor_s1_chipselect),       //                                              .chipselect
		.gpio_s1_address                                     (mm_interconnect_1_gpio_s1_address),              //                                       gpio_s1.address
		.gpio_s1_write                                       (mm_interconnect_1_gpio_s1_write),                //                                              .write
		.gpio_s1_readdata                                    (mm_interconnect_1_gpio_s1_readdata),             //                                              .readdata
		.gpio_s1_writedata                                   (mm_interconnect_1_gpio_s1_writedata),            //                                              .writedata
		.gpio_s1_chipselect                                  (mm_interconnect_1_gpio_s1_chipselect),           //                                              .chipselect
		.sysid_control_slave_address                         (mm_interconnect_1_sysid_control_slave_address),  //                           sysid_control_slave.address
		.sysid_control_slave_readdata                        (mm_interconnect_1_sysid_control_slave_readdata), //                                              .readdata
		.systimer_s1_address                                 (mm_interconnect_1_systimer_s1_address),          //                                   systimer_s1.address
		.systimer_s1_write                                   (mm_interconnect_1_systimer_s1_write),            //                                              .write
		.systimer_s1_readdata                                (mm_interconnect_1_systimer_s1_readdata),         //                                              .readdata
		.systimer_s1_writedata                               (mm_interconnect_1_systimer_s1_writedata),        //                                              .writedata
		.systimer_s1_chipselect                              (mm_interconnect_1_systimer_s1_chipselect),       //                                              .chipselect
		.sysuart_s1_address                                  (mm_interconnect_1_sysuart_s1_address),           //                                    sysuart_s1.address
		.sysuart_s1_write                                    (mm_interconnect_1_sysuart_s1_write),             //                                              .write
		.sysuart_s1_read                                     (mm_interconnect_1_sysuart_s1_read),              //                                              .read
		.sysuart_s1_readdata                                 (mm_interconnect_1_sysuart_s1_readdata),          //                                              .readdata
		.sysuart_s1_writedata                                (mm_interconnect_1_sysuart_s1_writedata),         //                                              .writedata
		.sysuart_s1_begintransfer                            (mm_interconnect_1_sysuart_s1_begintransfer),     //                                              .begintransfer
		.sysuart_s1_chipselect                               (mm_interconnect_1_sysuart_s1_chipselect),        //                                              .chipselect
		.vga_csr_address                                     (mm_interconnect_1_vga_csr_address),              //                                       vga_csr.address
		.vga_csr_write                                       (mm_interconnect_1_vga_csr_write),                //                                              .write
		.vga_csr_read                                        (mm_interconnect_1_vga_csr_read),                 //                                              .read
		.vga_csr_readdata                                    (mm_interconnect_1_vga_csr_readdata),             //                                              .readdata
		.vga_csr_writedata                                   (mm_interconnect_1_vga_csr_writedata)             //                                              .writedata
	);

	c4e_pcmplay_core_irq_mapper irq_mapper (
		.clk           (clk_100m_clk),                       //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),           // receiver4.irq
		.sender_irq    (nios2_tiny_irq_irq)                  //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (clk_25m_clk),                        //       receiver_clk.clk
		.sender_clk     (clk_100m_clk),                       //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver0_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_001 (
		.receiver_clk   (clk_25m_clk),                        //       receiver_clk.clk
		.sender_clk     (clk_100m_clk),                       //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_001_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver2_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_002 (
		.receiver_clk   (clk_25m_clk),                        //       receiver_clk.clk
		.sender_clk     (clk_100m_clk),                       //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_001_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_002_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver3_irq)            //             sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (clk_25m_clk),                    //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_tiny_debug_reset_request_reset),   // reset_in1.reset
		.clk            (clk_100m_clk),                           //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_100m_clk),                       //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_100m_clk),                       //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
